module top_module (
	input a,
	input b,
	input c,
	output w,
	output x,
	output y,
	output z  );
	
	assign w = a;
  assign y = b;
	assign x = b;
  assign z = c;

	
	
endmodule
